`define OP_ADD  'b00000
`define OP_SUB  'b00001

`define OP_SLL  'b00010
`define OP_SRL  'b00011
`define OP_SLA  'b00110
`define OP_SRA  'b00111

`define OP_SLT  'b00100
`define OP_SLTU 'b00101

`define OP_XOR  'b01000
`define OP_OR   'b01001
`define OP_AND  'b01010