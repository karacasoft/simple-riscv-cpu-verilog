`include "cpu_tests/test_common.vh"
`include "cpu.vh"

`define TEST_BRANCH(TNUM, RS2, RS1, RS2_VAL, RS1_VAL, OFFSET, INITIAL_PC, EXPECTED_PC, FUNCT3) `TEST_NUM(TNUM); \
    `RESET; \
    `REGISTER(RS1) = RS1_VAL; \
    `REGISTER(RS2) = RS2_VAL; \
    `PC = INITIAL_PC; \
    `SET_B_TYPE(OFFSET, RS2, RS1, FUNCT3, `BRANCH); \
    `DELAY_CYCLES(3); \
    `ASSERT_EQ(`PC, EXPECTED_PC); \

`define TEST_BEQ(TNUM, RS2, RS1, RS2_VAL, RS1_VAL, OFFSET, INITIAL_PC, EXPECTED_PC) `TEST_BRANCH(TNUM, RS2, RS1, RS2_VAL, RS1_VAL, OFFSET, INITIAL_PC, EXPECTED_PC, `FUNCT3_BEQ)
`define TEST_BNE(TNUM, RS2, RS1, RS2_VAL, RS1_VAL, OFFSET, INITIAL_PC, EXPECTED_PC) `TEST_BRANCH(TNUM, RS2, RS1, RS2_VAL, RS1_VAL, OFFSET, INITIAL_PC, EXPECTED_PC, `FUNCT3_BNE)
`define TEST_BLT(TNUM, RS2, RS1, RS2_VAL, RS1_VAL, OFFSET, INITIAL_PC, EXPECTED_PC) `TEST_BRANCH(TNUM, RS2, RS1, RS2_VAL, RS1_VAL, OFFSET, INITIAL_PC, EXPECTED_PC, `FUNCT3_BLT)
`define TEST_BGT(TNUM, RS2, RS1, RS2_VAL, RS1_VAL, OFFSET, INITIAL_PC, EXPECTED_PC) `TEST_BRANCH(TNUM, RS2, RS1, RS2_VAL, RS1_VAL, OFFSET, INITIAL_PC, EXPECTED_PC, `FUNCT3_BGT)
`define TEST_BLTU(TNUM, RS2, RS1, RS2_VAL, RS1_VAL, OFFSET, INITIAL_PC, EXPECTED_PC) `TEST_BRANCH(TNUM, RS2, RS1, RS2_VAL, RS1_VAL, OFFSET, INITIAL_PC, EXPECTED_PC, `FUNCT3_BLTU)
`define TEST_BGTU(TNUM, RS2, RS1, RS2_VAL, RS1_VAL, OFFSET, INITIAL_PC, EXPECTED_PC) `TEST_BRANCH(TNUM, RS2, RS1, RS2_VAL, RS1_VAL, OFFSET, INITIAL_PC, EXPECTED_PC, `FUNCT3_BGTU)