`define LSU_OP_SIZE_BYTE      2'b00
`define LSU_OP_SIZE_HALF_WORD 2'b01
`define LSU_OP_SIZE_WORD      2'b10

`define LSU_OP_UNSIGNED       1
`define LSU_OP_SIGNED         0